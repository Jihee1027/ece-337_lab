`timescale 1ns / 10ps

module adder_6bit #()();

endmodule

