`timescale 1ns / 10ps

module edge_rise(
  input logic clk, n_rst, async_in,
  output logic sync_out, edge_flag
);
  // Test default parameter values
  edge_det rise (.*);
  
endmodule
