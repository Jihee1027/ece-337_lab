`timescale 1ns / 10ps

module fsm ();


endmodule

