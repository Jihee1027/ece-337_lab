`timescale 1ns / 10ps

module rcu ();


endmodule

