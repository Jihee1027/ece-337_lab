`timescale 1ns / 10ps

module stp_4bit ();


endmodule

