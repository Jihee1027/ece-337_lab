`timescale 1ns / 10ps

module adder_128bit ();


endmodule

