`timescale 1ns / 10ps

module full_adder #()();

endmodule

