`timescale 1ns / 10ps

module rcv_block ();


endmodule

