`timescale 1ns / 10ps

module flex_counter #() ();


endmodule

